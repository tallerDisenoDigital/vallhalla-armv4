module RotationRightExtended #(parameter bus = 32)
	(input logic [bus-1:0] a, b,output logic [bus-1:0] s);
	//not implemented yet
	assign s = a;
	
endmodule
